magic
tech sky130A
magscale 1 2
timestamp 1605771998
<< nwell >>
rect -89 -36 119 236
<< nmos >>
rect 0 -366 30 -236
<< pmos >>
rect 0 0 30 200
<< ndiff >>
rect -53 -248 0 -236
rect -53 -354 -45 -248
rect -11 -354 0 -248
rect -53 -366 0 -354
rect 30 -248 84 -236
rect 30 -354 41 -248
rect 75 -354 84 -248
rect 30 -366 84 -354
<< pdiff >>
rect -53 184 0 200
rect -53 16 -45 184
rect -11 16 0 184
rect -53 0 0 16
rect 30 184 83 200
rect 30 16 41 184
rect 75 16 83 184
rect 30 0 83 16
<< ndiffc >>
rect -45 -354 -11 -248
rect 41 -354 75 -248
<< pdiffc >>
rect -45 16 -11 184
rect 41 16 75 184
<< poly >>
rect 0 200 30 226
rect 0 -37 30 0
rect -2 -39 32 -37
rect -18 -49 48 -39
rect -18 -83 -2 -49
rect 32 -83 48 -49
rect -18 -93 48 -83
rect -18 -149 48 -139
rect -18 -183 -2 -149
rect 32 -183 48 -149
rect -18 -193 48 -183
rect 0 -236 30 -193
rect 0 -392 30 -366
<< polycont >>
rect -2 -83 32 -49
rect -2 -183 32 -149
<< locali >>
rect -70 184 -11 200
rect -70 16 -45 184
rect -70 0 -11 16
rect 41 184 100 200
rect 75 16 100 184
rect 41 0 100 16
rect -70 -232 -36 0
rect -2 -49 32 -33
rect -2 -99 32 -83
rect -2 -149 32 -133
rect -2 -199 32 -183
rect 66 -232 100 0
rect -70 -248 -11 -232
rect -70 -354 -45 -248
rect -70 -370 -11 -354
rect 41 -248 100 -232
rect 75 -354 100 -248
rect 41 -370 100 -354
<< labels >>
rlabel polycont -2 -83 32 -49 1 Cnot
port 2 n
rlabel polycont -2 -183 32 -149 1 C
port 1 n
rlabel locali -70 -248 -36 16 1 A
port 3 n
rlabel locali 66 -248 100 16 1 B
port 4 n
<< end >>

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO transmission_gate_cell
  CLASS CORE ;
  FOREIGN transmission_gate_cell ;
  ORIGIN 0.470 1.970 ;
  SIZE 1.090 BY 3.200 ;
  SITE unithd ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.097500 ;
    PORT
      LAYER li1 ;
        RECT -0.010 -0.995 0.160 -0.665 ;
    END
  END C
  PIN Cnot
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.150000 ;
    PORT
      LAYER li1 ;
        RECT -0.010 -0.495 0.160 -0.165 ;
    END
  END Cnot
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.437250 ;
    PORT
      LAYER li1 ;
        RECT -0.350 0.000 -0.055 1.000 ;
        RECT -0.350 -1.160 -0.180 0.000 ;
        RECT -0.350 -1.850 -0.055 -1.160 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440500 ;
    PORT
      LAYER li1 ;
        RECT 0.205 0.000 0.500 1.000 ;
        RECT 0.330 -1.160 0.500 0.000 ;
        RECT 0.205 -1.850 0.500 -1.160 ;
    END
  END B
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT -0.470 0.750 0.620 1.230 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT -0.470 -1.970 0.620 -1.490 ;
    END
  END VGND
END transmission_gate_cell
END LIBRARY


(* blackbox *)
module transmission_gate_cell(inout a, inout b, input c, input c_not);
endmodule

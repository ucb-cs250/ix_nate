(* blackbox *)
module transmission_gate(inout a, inout b, input c, input c_not);
endmodule

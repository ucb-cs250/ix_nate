magic
tech sky130A
magscale 1 2
timestamp 1606263321
<< nwell >>
rect -38 261 315 584
<< pwell >>
rect 11 -19 45 15
<< scnmos >>
rect 165 47 195 177
<< pmoshvt >>
rect 81 297 111 497
<< ndiff >>
rect 29 161 165 177
rect 29 67 37 161
rect 71 148 165 161
rect 71 67 121 148
rect 155 67 165 148
rect 29 47 165 67
rect 195 159 247 177
rect 195 64 205 159
rect 239 64 247 159
rect 195 47 247 64
<< pdiff >>
rect 29 480 81 497
rect 29 383 37 480
rect 71 383 81 480
rect 29 349 81 383
rect 29 315 37 349
rect 71 315 81 349
rect 29 297 81 315
rect 111 477 247 497
rect 111 325 121 477
rect 155 383 205 477
rect 239 383 247 477
rect 155 349 247 383
rect 155 325 205 349
rect 111 315 205 325
rect 239 315 247 349
rect 111 297 247 315
<< ndiffc >>
rect 37 67 71 161
rect 121 67 155 148
rect 205 64 239 159
<< pdiffc >>
rect 37 383 71 480
rect 37 315 71 349
rect 121 325 155 477
rect 205 383 239 477
rect 205 315 239 349
<< poly >>
rect 81 497 111 523
rect 81 265 111 297
rect 51 249 117 265
rect 51 215 67 249
rect 101 215 117 249
rect 51 199 117 215
rect 159 259 225 275
rect 159 225 175 259
rect 209 225 225 259
rect 159 209 225 225
rect 165 177 195 209
rect 165 21 195 47
<< polycont >>
rect 67 215 101 249
rect 175 225 209 259
<< locali >>
rect 9 495 71 496
rect -5 480 71 495
rect -5 383 37 480
rect -5 349 71 383
rect -5 315 37 349
rect -5 299 71 315
rect 112 477 277 493
rect 112 325 121 477
rect 155 383 205 477
rect 239 383 277 477
rect 155 349 277 383
rect 155 325 205 349
rect 112 315 205 325
rect 239 315 277 349
rect 112 309 277 315
rect -5 164 33 299
rect 67 249 101 265
rect 67 199 101 215
rect 175 259 209 275
rect 175 209 209 225
rect 243 175 277 309
rect -5 161 164 164
rect -5 67 37 161
rect 71 148 164 161
rect 71 67 121 148
rect 155 67 164 148
rect -5 51 164 67
rect 205 159 277 175
rect 239 64 277 159
rect 205 49 277 64
rect 205 48 276 49
<< metal1 >>
rect 0 496 276 592
rect 0 -48 276 48
<< labels >>
rlabel nwell s 11 -19 45 15 1 VNB
rlabel metal1 0 -48 276 48 1 VGND
port 1 n ground bidirectional abutment
rlabel metal1 18 530 52 564 1 VPB
rlabel metal1 0 496 276 592 1 VPWR
port 2 n ground bidirectional abutment
rlabel locali -5 51 33 495 1 A
port 3 n signal bidirectional
rlabel locali 243 49 277 493 1 B
port 4 n signal bidirectional
rlabel polycont 67 215 101 249 1 Cnot
port 5 n signal input
rlabel polycont 175 225 209 259 1 C
port 6 n signal input
<< properties >>
string LEFclass CORE
string LEFsite unithd
string FIXED_BBOX -5 0 282 544
string LEFsymmetry X Y R90
string LEFsource user
<< end >>

(* blackbox *)
module transmission_gate(inout a, inout b, input c);
endmodule

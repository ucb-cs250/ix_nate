(* blackbox *)
module transmission_gate_cell(inout A, inout B, input C, input Cnot);
endmodule

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO transmission_gate_cell
  CLASS CORE ;
  FOREIGN transmission_gate_cell ;
  ORIGIN 0.025 0.000 ;
  SIZE 1.435 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.702000 ;
    PORT
      LAYER li1 ;
        RECT 0.045 2.475 0.355 2.480 ;
        RECT -0.025 1.495 0.355 2.475 ;
        RECT -0.025 0.820 0.165 1.495 ;
        RECT -0.025 0.255 0.820 0.820 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.849000 ;
    PORT
      LAYER li1 ;
        RECT 0.560 1.545 1.385 2.465 ;
        RECT 1.215 0.875 1.385 1.545 ;
        RECT 1.025 0.245 1.385 0.875 ;
        RECT 1.025 0.240 1.380 0.245 ;
    END
  END B
  PIN Cnot
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.150000 ;
    PORT
      LAYER li1 ;
        RECT 0.335 0.995 0.505 1.325 ;
    END
  END Cnot
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.097500 ;
    PORT
      LAYER li1 ;
        RECT 0.875 1.045 1.045 1.375 ;
    END
  END C
END transmission_gate_cell
END LIBRARY


* SPICE3 file created from /home/nate/Projects/cs250/ix_nate/transgate.ext - technology: sky130A

.option scale=5000u

X0 B C A $SUB sky130_fd_pr__nfet_01v8 w=50 l=30
X1 B Cnot A w_n68_58# sky130_fd_pr__pfet_01v8 w=54 l=30

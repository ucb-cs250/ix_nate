VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO transmission_gate_cell
  CLASS CORE ;
  FOREIGN transmission_gate_cell ;
  ORIGIN 0.110 0.000 ;
  SIZE 1.580 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN Cnot
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.150000 ;
    PORT
      LAYER li1 ;
        RECT 0.335 0.995 0.505 1.325 ;
    END
  END Cnot
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.097500 ;
    PORT
      LAYER li1 ;
        RECT 0.875 1.000 1.045 1.330 ;
    END
  END C
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.712000 ;
    PORT
      LAYER li1 ;
        RECT -0.025 1.495 0.355 2.465 ;
        RECT -0.025 0.820 0.165 1.495 ;
        RECT -0.025 0.255 0.820 0.820 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.852250 ;
    PORT
      LAYER li1 ;
        RECT 0.560 1.545 1.385 2.465 ;
        RECT 1.215 0.830 1.385 1.545 ;
        RECT 0.995 0.255 1.385 0.830 ;
    END
  END B
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT -0.110 2.480 1.470 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT -0.110 -0.240 1.470 0.240 ;
    END
  END VGND
END transmission_gate_cell
END LIBRARY


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO transmission_gate
  CLASS BLOCK ;
  FOREIGN transmission_gate ;
  ORIGIN 0.340 0.730 ;
  SIZE 1.090 BY 2.000 ;
  PIN B
    ANTENNADIFFAREA 0.150800 ;
    PORT
      LAYER li1 ;
        RECT 0.320 -0.340 0.530 0.830 ;
    END
  END B
  PIN A
    ANTENNADIFFAREA 0.150800 ;
    PORT
      LAYER li1 ;
        RECT -0.120 -0.340 0.090 0.830 ;
    END
  END A
  PIN Cnot
    ANTENNAGATEAREA 0.040500 ;
    PORT
      LAYER li1 ;
        RECT 0.040 1.050 0.370 1.220 ;
    END
  END Cnot
  PIN C
    ANTENNAGATEAREA 0.037500 ;
    PORT
      LAYER li1 ;
        RECT 0.040 -0.680 0.370 -0.510 ;
    END
  END C
END transmission_gate
END LIBRARY

